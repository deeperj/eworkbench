** Profile: "FULLADD-SWEEP"  [ E:\OrCAD\16.2\kits\postbeta\uploadedkits\October5\orcadFlowTutDoc\doc\flowtut\tutorial_example\Flowtut\partial\fulladd-PSpiceFiles\FULLADD\SWEEP.sim ] 

** Creating circuit file "SWEEP.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.STMLIB "../../../fulladd-pspicefiles/fulladd/sweep/input.stl" 
* From [PSPICE NETLIST] section of E:\OrCAD\OrCAD_16.2\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 100us 0 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\FULLADD.net" 


.END
